module or1(input a, input b, output c);
assign c= a | b;
endmodule
